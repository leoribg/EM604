library verilog;
use verilog.vl_types.all;
entity project2_vlg_vec_tst is
end project2_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity project2_TB is
end project2_TB;

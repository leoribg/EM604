library verilog;
use verilog.vl_types.all;
entity divisorSM_vlg_vec_tst is
end divisorSM_vlg_vec_tst;

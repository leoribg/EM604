library verilog;
use verilog.vl_types.all;
entity projeto_vlg_vec_tst is
end projeto_vlg_vec_tst;
